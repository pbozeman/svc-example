`include "svc.sv"

`include "svc_soc_sim.sv"

//
// Standalone interactive simulation for RISC-V bubble sort demo
//
// Architecture-generic: hex file path set by Makefile via RV_BUBBLE_SORT_HEX define
//
// Usage:
//   make sw
//   make rv_bubble_sort_i_sim        # RV32I variant
//   make rv_bubble_sort_im_sim       # RV32IM variant
//   make rv_bubble_sort_i_zmmul_sim  # RV32I_Zmmul variant (hardware multiply)
//
module rv_bubble_sort_sim;
  //
  // Shared configuration from Makefile defines
  //
  `include "rv_sim_config.svh"

  //
  // Program-specific configuration
  //
  localparam int WATCHDOG_CYCLES = 500_000;  // 20ms at 25MHz

  //
  // SOC simulation with CPU, peripherals, and lifecycle management
  //
  svc_soc_sim #(
      // Clock and timing
      .CLOCK_FREQ_MHZ (25),
      .WATCHDOG_CYCLES(WATCHDOG_CYCLES),
      // Memory configuration
      .IMEM_DEPTH     (IMEM_DEPTH),
      .DMEM_DEPTH     (DMEM_DEPTH),
      .IMEM_INIT      (MEM_INIT),
      .DMEM_INIT      (MEM_INIT),
      // CPU architecture (from rv_sim_config.svh)
      .MEM_TYPE       (MEM_TYPE),
      .PIPELINED      (PIPELINED),
      .FWD_REGFILE    (FWD_REGFILE),
      .FWD            (FWD),
      .BPRED          (BPRED),
      .BTB_ENABLE     (BTB_ENABLE),
      .EXT_ZMMUL      (EXT_ZMMUL),
      .EXT_M          (EXT_M),
      // Peripherals
      .BAUD_RATE      (115_200),
      // Debug/reporting
      .PREFIX         ("bubble"),
      .SW_PATH        ("sw/bubble_sort/main.c")
  ) sim ();

  //
  // Optional: Generate VCD for waveform viewing
  //
  // initial begin
  //   $dumpfile("rv_bubble_sort_sim.vcd");
  //   $dumpvars(0, rv_bubble_sort_sim);
  // end

endmodule
